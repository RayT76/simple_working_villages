5:local _={};_[1]="default:gravel";_[2]="default:wood";_[3]="inventory";_[4]="default:fence_wood";_[5]="default:torch_wall";_[6]="default:dirt";_[7]="default:ladder_wood";return {{x=0,y=1,param1=14,z=0,name=_[4]},{x=0,y=1,param1=15,z=1,name=_[4]},{x=0,y=1,param1=15,z=2,name=_[4]},{x=0,y=1,param1=15,z=3,name=_[4]},{x=0,y=1,param1=15,z=4,name=_[4]},{x=0,y=1,param1=31,z=5,name=_[4]},{x=0,y=1,param1=47,z=6,name=_[4]},{x=0,y=1,param1=63,z=7,name=_[4]},{x=0,y=1,param1=79,z=8,name=_[4]},{x=0,y=1,param1=63,z=9,name=_[4]},{x=0,y=1,param1=47,z=10,name=_[4]},{x=0,y=1,param1=63,z=11,name=_[4]},{x=0,y=1,param1=79,z=12,name=_[4]},{x=0,y=1,param1=95,z=13,name=_[4]},{x=0,y=1,param1=79,z=14,name=_[4]},{x=0,y=1,param1=63,z=15,name=_[4]},{x=0,y=1,param1=47,z=16,name=_[4]},{x=0,y=1,param1=31,z=17,name=_[4]},{x=0,y=1,param1=15,z=18,name=_[4]},{x=0,y=1,param1=15,z=19,name=_[4]},{x=0,y=2,z=0,name=_[6]},{x=0,y=3,z=0,name=_[6]},{x=1,y=1,param1=15,z=0,name=_[4]},{x=1,y=1,param1=15,z=19,name=_[4]},{x=2,y=1,param1=15,z=0,name=_[4]},{x=2,y=1,param1=15,z=19,name=_[4]},{x=3,y=1,param1=15,z=0,name=_[4]},{x=3,y=1,param1=15,z=19,name=_[4]},{x=4,y=1,param1=15,z=0,name=_[4]},{x=4,y=1,param1=31,z=19,name=_[4]},{x=5,y=1,param1=31,z=0,name=_[4]},{x=5,y=1,z=7,name=_[2]},{x=5,y=1,z=8,name=_[2]},{x=5,y=1,z=9,name=_[2]},{x=5,y=1,z=10,name=_[2]},{x=5,y=1,z=11,name=_[2]},{x=5,y=1,z=12,name=_[2]},{x=5,y=1,param1=47,z=19,name=_[4]},{x=5,y=2,param1=158,z=7,name=_[4]},{x=5,y=2,param1=174,z=8,name=_[4]},{x=5,y=2,param1=158,z=9,name=_[4]},{x=5,y=2,param1=142,z=10,name=_[4]},{x=5,y=2,param1=158,z=11,name=_[4]},{x=5,y=2,param1=142,z=12,name=_[4]},{x=5,y=3,z=7,name=_[2]},{x=5,y=3,z=8,name=_[2]},{x=5,y=3,z=9,name=_[2]},{x=5,y=3,z=10,name=_[2]},{x=5,y=3,z=11,name=_[2]},{x=5,y=3,z=12,name=_[2]},{x=5,y=4,z=7,name=_[2]},{x=5,y=4,z=8,name=_[2]},{x=5,y=4,z=9,name=_[2]},{x=5,y=4,z=10,name=_[2]},{x=5,y=4,z=11,name=_[2]},{x=5,y=4,z=12,name=_[2]},{x=6,y=0,z=8,name=_[1]},{x=6,y=0,z=9,name=_[1]},{x=6,y=0,z=10,name=_[1]},{x=6,y=0,z=11,name=_[1]},{x=6,y=1,param1=47,z=0,name=_[4]},{x=6,y=1,z=7,name=_[2]},{x=6,meta={fields={infotext="\27(T@default)Chest\27E"},[_[3]]={main={"","","","","","","","","","","","","","","","","","","","","","","","","","","","","","","",""}}},param2=2,y=1,param1=174,z=8,name="default:chest"},{x=6,y=1,z=12,name=_[2]},{x=6,y=1,param1=63,z=19,name=_[4]},{x=6,y=2,param1=174,z=7,name=_[4]},{x=6,y=2,z=12,name=_[2]},{x=6,y=3,z=7,name=_[2]},{x=6,param2=5,y=3,param1=206,z=8,name=_[5]},{x=6,y=3,z=12,name=_[2]},{x=6,y=4,z=7,name=_[2]},{x=6,y=4,z=8,name=_[2]},{x=6,y=4,z=9,name=_[2]},{x=6,y=4,z=10,name=_[2]},{x=6,y=4,z=11,name=_[2]},{x=6,y=4,z=12,name=_[2]},{x=7,y=0,z=8,name=_[1]},{x=7,y=0,z=9,name=_[1]},{x=7,y=0,z=10,name=_[1]},{x=7,y=0,z=11,name=_[1]},{x=7,y=0,z=12,name=_[1]},{x=7,y=0,z=13,name=_[1]},{x=7,y=0,z=14,name=_[1]},{x=7,y=0,z=15,name=_[1]},{x=7,y=0,z=16,name=_[1]},{x=7,y=0,z=17,name=_[1]},{x=7,y=0,z=18,name=_[1]},{x=7,y=0,z=19,name=_[1]},{x=7,y=1,param1=31,z=0,name=_[4]},{x=7,y=1,z=7,name=_[2]},{x=7,param2=5,y=1,param1=159,z=8,name=_[7]},{x=7,meta={fields={state="1"},[_[3]]={}},param2=3,y=1,param1=158,z=12,name="doors:door_wood_c"},{x=7,y=2,z=7,name=_[2]},{x=7,param2=5,y=2,param1=175,z=8,name=_[7]},{x=7,param2=2,y=2,param1=174,z=12,name="doors:hidden"},{x=7,y=3,z=7,name=_[2]},{x=7,param2=5,y=3,param1=191,z=8,name=_[7]},{x=7,param2=4,y=3,param1=204,z=11,name=_[5]},{x=7,y=3,z=12,name=_[2]},{x=7,param2=5,y=3,param1=207,z=13,name=_[5]},{x=7,y=4,z=7,name=_[2]},{x=7,param2=5,y=4,param1=175,z=8,name=_[7]},{x=7,y=4,z=9,name=_[2]},{x=7,y=4,z=10,name=_[2]},{x=7,y=4,z=11,name=_[2]},{x=7,y=4,z=12,name=_[2]},{x=8,y=0,z=8,name=_[1]},{x=8,y=0,z=9,name=_[1]},{x=8,y=0,z=10,name=_[1]},{x=8,y=0,z=11,name=_[1]},{x=8,y=1,param1=15,z=0,name=_[4]},{x=8,y=1,z=7,name=_[2]},{x=8,param2=2,y=1,param1=142,z=8,name="beds:bed_top"},{x=8,param2=2,y=1,param1=125,z=9,name="beds:bed_bottom"},{x=8,y=1,z=12,name=_[2]},{x=8,y=1,param1=63,z=19,name=_[4]},{x=8,y=2,param1=142,z=7,name=_[4]},{x=8,y=2,z=12,name=_[2]},{x=8,y=3,z=7,name=_[2]},{x=8,y=3,z=12,name=_[2]},{x=8,y=4,z=7,name=_[2]},{x=8,y=4,z=8,name=_[2]},{x=8,y=4,z=9,name=_[2]},{x=8,y=4,z=10,name=_[2]},{x=8,y=4,z=11,name=_[2]},{x=8,y=4,z=12,name=_[2]},{x=9,y=1,param1=15,z=0,name=_[4]},{x=9,y=1,z=7,name=_[2]},{x=9,y=1,z=8,name=_[2]},{x=9,y=1,z=9,name=_[2]},{x=9,y=1,z=10,name=_[2]},{x=9,y=1,z=11,name=_[2]},{x=9,y=1,z=12,name=_[2]},{x=9,y=1,param1=47,z=19,name=_[4]},{x=9,y=2,param1=126,z=7,name=_[4]},{x=9,y=2,param1=142,z=8,name=_[4]},{x=9,y=2,param1=126,z=9,name=_[4]},{x=9,y=2,param1=142,z=10,name=_[4]},{x=9,y=2,param1=158,z=11,name=_[4]},{x=9,y=2,param1=142,z=12,name=_[4]},{x=9,y=3,z=7,name=_[2]},{x=9,y=3,z=8,name=_[2]},{x=9,y=3,z=9,name=_[2]},{x=9,y=3,z=10,name=_[2]},{x=9,y=3,z=11,name=_[2]},{x=9,y=3,z=12,name=_[2]},{x=9,y=4,z=7,name=_[2]},{x=9,y=4,z=8,name=_[2]},{x=9,y=4,z=9,name=_[2]},{x=9,y=4,z=10,name=_[2]},{x=9,y=4,z=11,name=_[2]},{x=9,y=4,z=12,name=_[2]},{x=10,y=1,param1=15,z=0,name=_[4]},{x=10,y=1,param1=31,z=19,name=_[4]},{x=11,y=1,param1=15,z=0,name=_[4]},{x=11,y=1,param1=15,z=19,name=_[4]},{x=12,y=1,param1=15,z=0,name=_[4]},{x=12,y=1,param1=15,z=19,name=_[4]},{x=13,y=1,param1=15,z=0,name=_[4]},{x=13,y=1,param1=31,z=19,name=_[4]},{x=14,y=1,param1=15,z=0,name=_[4]},{x=14,y=1,param1=15,z=1,name=_[4]},{x=14,y=1,param1=15,z=2,name=_[4]},{x=14,y=1,param1=15,z=3,name=_[4]},{x=14,y=1,param1=15,z=4,name=_[4]},{x=14,y=1,param1=15,z=5,name=_[4]},{x=14,y=1,param1=15,z=6,name=_[4]},{x=14,y=1,param1=31,z=7,name=_[4]},{x=14,y=1,param1=47,z=8,name=_[4]},{x=14,y=1,param1=31,z=9,name=_[4]},{x=14,y=1,param1=47,z=10,name=_[4]},{x=14,y=1,param1=63,z=11,name=_[4]},{x=14,y=1,param1=47,z=12,name=_[4]},{x=14,y=1,param1=63,z=13,name=_[4]},{x=14,y=1,param1=63,z=14,name=_[4]},{x=14,y=1,param1=47,z=15,name=_[4]},{x=14,y=1,param1=31,z=16,name=_[4]},{x=14,y=1,param1=15,z=17,name=_[4]},{x=14,y=1,param1=31,z=18,name=_[4]},{x=14,y=1,param1=47,z=19,name=_[4]}}