5:local _={};_[1]="default:fence_wood";_[2]="homedecor:kitchen_chair_wood";_[3]="beds:bed_bottom";_[4]="default:chest";_[5]="default:torch";_[6]="infotext";_[7]="\27(T@default)Chest\27E";_[8]="beds:bed_top";_[9]="inventory";return {{x=0,y=0,param1=191,z=0,name=_[1]},{x=0,y=0,param1=175,z=1,name=_[1]},{x=0,y=0,param1=159,z=2,name=_[1]},{x=0,y=0,param1=143,z=3,name=_[1]},{x=0,y=0,param1=143,z=5,name=_[1]},{x=0,y=0,param1=159,z=6,name=_[1]},{x=0,y=0,param1=175,z=7,name=_[1]},{x=0,y=0,param1=191,z=8,name=_[1]},{x=0,param2=1,y=1,param1=207,z=0,name=_[5]},{x=0,param2=1,y=1,param1=207,z=8,name=_[5]},{x=1,y=0,param1=175,z=0,name=_[1]},{x=1,y=0,param1=175,z=8,name=_[1]},{x=2,y=0,param1=159,z=0,name=_[1]},{x=2,y=0,param1=159,z=8,name=_[1]},{x=3,y=0,param1=143,z=0,name=_[1]},{x=3,y=0,param1=143,z=8,name=_[1]},{x=5,y=0,param1=111,z=0,name=_[1]},{x=5,y=0,param1=111,z=8,name=_[1]},{x=6,y=0,param1=127,z=0,name=_[1]},{x=6,y=0,param1=95,z=8,name=_[1]},{x=7,y=0,param1=143,z=0,name=_[1]},{x=7,y=0,param1=79,z=8,name=_[1]},{x=8,y=0,param1=159,z=0,name=_[1]},{x=8,y=0,param1=175,z=1,name=_[1]},{x=8,y=0,param1=191,z=2,name=_[1]},{x=8,y=0,param1=175,z=3,name=_[1]},{x=8,y=0,param1=143,z=5,name=_[1]},{x=8,y=0,param1=127,z=6,name=_[1]},{x=8,y=0,param1=111,z=7,name=_[1]},{x=8,y=0,param1=95,z=8,name=_[1]},{x=9,y=0,param1=175,z=0,name=_[1]},{x=9,y=0,param1=142,z=6,name=_[3]},{x=9,y=0,param1=126,z=7,name=_[8]},{x=9,y=0,param1=111,z=8,name=_[1]},{x=10,y=0,param1=191,z=0,name=_[1]},{x=10,meta={fields={layer_2="20",layer_3="21",layer_1="19"},[_[9]]={}},param2=2,y=0,param1=223,z=2,name="fake_fire:fancy_fire"},{x=10,y=0,param1=127,z=8,name=_[1]},{x=11,y=0,param1=175,z=0,name=_[1]},{x=11,param2=5,y=0,param1=126,z=7,name=_[2]},{x=11,y=0,param1=111,z=8,name=_[1]},{x=12,y=0,param1=159,z=0,name=_[1]},{x=12,y=0,param1=110,z=7,name="homedecor:table"},{x=12,y=0,param1=127,z=8,name=_[1]},{x=13,y=0,param1=143,z=0,name=_[1]},{x=13,param2=1,y=0,param1=158,z=1,name=_[3]},{x=13,param2=4,y=0,param1=126,z=7,name=_[2]},{x=13,y=0,param1=143,z=8,name=_[1]},{x=14,y=0,param1=159,z=0,name=_[1]},{x=14,param2=1,y=0,param1=142,z=1,name=_[8]},{x=14,y=0,param1=159,z=8,name=_[1]},{x=15,y=0,param1=175,z=0,name=_[1]},{x=15,meta={fields={[_[6]]=_[7]},[_[9]]={main={"","","","","","","","","","","","","","","","","","","","","","","","","","","","","","","",""}}},param2=2,y=0,param1=158,z=1,name=_[4]},{x=15,meta={fields={[_[6]]=_[7]},[_[9]]={main={"","","","","","","","","","","","","","","","","","","","","","","","","","","","","","","",""}}},y=0,param1=158,z=7,name=_[4]},{x=15,y=0,param1=175,z=8,name=_[1]},{x=16,y=0,param1=191,z=0,name=_[1]},{x=16,y=0,param1=175,z=1,name=_[1]},{x=16,y=0,param1=159,z=2,name=_[1]},{x=16,y=0,param1=143,z=3,name=_[1]},{x=16,y=0,param1=143,z=5,name=_[1]},{x=16,y=0,param1=159,z=6,name=_[1]},{x=16,y=0,param1=175,z=7,name=_[1]},{x=16,y=0,param1=191,z=8,name=_[1]},{x=16,param2=1,y=1,param1=207,z=0,name=_[5]},{x=16,param2=1,y=1,param1=207,z=8,name=_[5]}}